`timescale 1ns / 1ps

module uart_test_top(
    input  wire       clk,          // ϵͳʱ�� (100MHz)
    input  wire       rst_n,        // ��λ�ź� (�͵�ƽ��Ч���ɰ󶨵�һ�������򿪹�)
    input  wire       uart_rx,      // UART ��������
    output wire       uart_tx,      // UART ��������
    output wire [7:0] led           // LED ��ʾ���յ�������
);

    // ==========================================
    // ��������
    // ==========================================
    parameter CLK_FREQ  = 100_000_000; // �������İ���ʵ��ʱ��Ƶ���޸�
    parameter BAUD_RATE = 115200;      // ������

    // ==========================================
    // �ڲ��ź�
    // ==========================================
    wire [7:0] rx_data;
    wire       rx_done;
    wire       tx_busy;
    
    reg  [7:0] tx_data_reg;
    reg        tx_start_reg;

    // �����յ�������ֱ�����ӵ� LED
    // ע�⣺����Ǹ��߼�LED���͵�ƽ������������Ҫȡ������ assign led = ~rx_data;
    assign led = rx_data; 

    // ==========================================
    // ģ������
    // ==========================================

    // 1. ���ڽ���ģ��
    uart_rx #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) u_rx (
        .clk(clk),
        .rst_n(~rst_n),
        .rx(uart_rx),
        .rx_data(rx_data),
        .rx_done(rx_done)
    );

    // 2. ���ڷ���ģ��
    uart_tx #(
        .CLK_FREQ(CLK_FREQ),
        .BAUD_RATE(BAUD_RATE)
    ) u_tx (
        .clk(clk),
        .rst_n(~rst_n),
        .tx_start(tx_start_reg),
        .tx_data(tx_data_reg),
        .tx(uart_tx),
        .tx_busy(tx_busy)
    );

    // ==========================================
    // �ػ��߼� (Loopback Logic)
    // ==========================================
    // �����յ����� (rx_done ����) ʱ��������Ͷ˲�æ���򴥷�����
    always @(posedge clk or posedge rst_n) begin
        if (rst_n) begin
            tx_start_reg <= 1'b0;
            tx_data_reg  <= 8'd0;
        end else begin
            // Ĭ�����������źţ�������ʽ��
            tx_start_reg <= 1'b0;

            // ��������ɣ��ҷ���ģ�����ʱ
            if (rx_done && !tx_busy) begin
                tx_data_reg  <= rx_data; // �����յ������ݸ����Ͷ�
                tx_start_reg <= 1'b1;    // ����һ��ʱ�����ڵĿ�ʼ����
            end
        end
    end

endmodule