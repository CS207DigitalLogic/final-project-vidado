`timescale 1ns / 1ps

module matrix_displayer(
    input wire clk,
    input wire rst_n,
    
    // �����ź�
    input wire start,           // ��ʼ��ʾ������
    output reg busy,            // ģ��æ�ź�
    
    // �����������
    input wire [2:0] matrix_row, // ��������
    input wire [2:0] matrix_col, // ��������
    
    // ���� Storage �� 25 ������
    input wire [7:0] d0,  input wire [7:0] d1,  input wire [7:0] d2,  input wire [7:0] d3,  input wire [7:0] d4,
    input wire [7:0] d5,  input wire [7:0] d6,  input wire [7:0] d7,  input wire [7:0] d8,  input wire [7:0] d9,
    input wire [7:0] d10, input wire [7:0] d11, input wire [7:0] d12, input wire [7:0] d13, input wire [7:0] d14,
    input wire [7:0] d15, input wire [7:0] d16, input wire [7:0] d17, input wire [7:0] d18, input wire [7:0] d19,
    input wire [7:0] d20, input wire [7:0] d21, input wire [7:0] d22, input wire [7:0] d23, input wire [7:0] d24,

    // UART TX �ӿ�
    output reg [7:0] tx_data,
    output reg       tx_start,
    input  wire      tx_busy
);

    // ״̬������
    localparam S_IDLE       = 0;
    localparam S_PREPARE    = 1; // ��������
    localparam S_SEND_DIGIT = 2; // ��������
    localparam S_WAIT_DIGIT = 3; // �ȴ����ַ���
    localparam S_SEND_SEP   = 4; // ���ͷָ���(�ո����)
    localparam S_WAIT_SEP   = 5; // �ȴ��ָ�������
    localparam S_DONE       = 6;

    reg [3:0] state;
    reg [2:0] r_cnt; // �м���
    reg [2:0] c_cnt; // �м���
    
    // �ڲ����ݻ��棨��ֹ��ʾ������ storage ���ˣ�
    reg [7:0] data_cache [24:0]; 
    reg [7:0] current_val;

    // ����ѡ���߼������� (r, c) ѡ����Ӧ������
    wire [4:0] current_index = r_cnt * matrix_col + c_cnt;

    // ����תASCII
    function [7:0] int2ascii;
        input [7:0] val;
        begin
            int2ascii = val + "0"; // �򵥴���0-9�����֧����λ����Ҫ�������߼�
        end
    endfunction

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_IDLE;
            busy <= 0;
            tx_start <= 0;
            tx_data <= 0;
            r_cnt <= 0;
            c_cnt <= 0;
        end else begin
            // Ĭ������ Start
            tx_start <= 0;

            case (state)
                S_IDLE: begin
                    busy <= 0;
                    if (start) begin
                        busy <= 1;
                        state <= S_PREPARE;
                    end
                end

                S_PREPARE: begin
                    // ������˿ڵ��������浽�ڲ����棬��֤��ʾʱ�����ȶ�
                    data_cache[0]<=d0;   data_cache[1]<=d1;   data_cache[2]<=d2;   data_cache[3]<=d3;   data_cache[4]<=d4;
                    data_cache[5]<=d5;   data_cache[6]<=d6;   data_cache[7]<=d7;   data_cache[8]<=d8;   data_cache[9]<=d9;
                    data_cache[10]<=d10; data_cache[11]<=d11; data_cache[12]<=d12; data_cache[13]<=d13; data_cache[14]<=d14;
                    data_cache[15]<=d15; data_cache[16]<=d16; data_cache[17]<=d17; data_cache[18]<=d18; data_cache[19]<=d19;
                    data_cache[20]<=d20; data_cache[21]<=d21; data_cache[22]<=d22; data_cache[23]<=d23; data_cache[24]<=d24;
                    
                    r_cnt <= 0;
                    c_cnt <= 0;
                    state <= S_SEND_DIGIT;
                end

                S_SEND_DIGIT: begin
                    if (!tx_busy) begin
                        // 1. ȡ����ǰ���ֲ�תASCII
                        current_val = data_cache[current_index];
                        tx_data <= int2ascii(current_val);
                        tx_start <= 1;
                        state <= S_WAIT_DIGIT;
                    end
                end

                S_WAIT_DIGIT: begin
                    // �ȴ�����æµ���������߷������
                    // һ������ֻҪ����start����һ����tx_busy�ͻ��ߣ��������ǿ��Լ򵥸�����ʱ
                    // ������ü򵥵�״̬��ת����Ϊ tx_busy �߼�ͨ����������Ӧ
                    state <= S_SEND_SEP;
                end

                S_SEND_SEP: begin
                    if (!tx_busy) begin
                        // �ж�����ĩ�����м�
                        if (c_cnt == matrix_col - 1) begin
                            tx_data <= 8'h0A; // ���� (Line Feed)
                            // ĳЩ�ն˿�����Ҫ 0D 0A�������Ϊ \n
                        end else begin
                            tx_data <= 8'h20; // �ո�
                        end
                        tx_start <= 1;
                        state <= S_WAIT_SEP;
                    end
                end

                S_WAIT_SEP: begin
                    if (!tx_busy) begin // �ȴ��ָ�������
                        // ���¼�����
                        if (c_cnt == matrix_col - 1) begin
                            c_cnt <= 0;
                            if (r_cnt == matrix_row - 1) begin
                                state <= S_DONE;
                            end else begin
                                r_cnt <= r_cnt + 1;
                                state <= S_SEND_DIGIT;
                            end
                        end else begin
                            c_cnt <= c_cnt + 1;
                            state <= S_SEND_DIGIT;
                        end
                    end
                end

                S_DONE: begin
                    busy <= 0;
                    state <= S_IDLE;
                end
            endcase
        end
    end

endmodule